module OwO;
  initial begin
    $display("OwO");
  end
endmodule
